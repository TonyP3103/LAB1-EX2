module wrapper ( 
						input logic [8:0] SW,
						input logic [1:0] KEY,
						output logic [9:0] LEDR,
						output logic [6:0] HEX0,HEX1,HEX2,HEX3);
						
ex2 wrapp (.clk(KEY[1]),.rst(KEY[0]),.a(SW),.out(LEDR[7:0]),.carry_out(LEDR[8]),.ovr(LEDR[9]),.c_in(SW[8]));

always_comb begin
case (SW[3:0])
	    4'b0000: HEX0 = 7'b1000000;//0
	    4'b0001: HEX0 = 7'b1111001;//1
	    4'b0010: HEX0 = 7'b0100100;//2
	    4'b0011: HEX0 = 7'b0110000;//3
	    4'b0100: HEX0 = 7'b0011001;//4
	    4'b0101: HEX0 = 7'b0010010;//5
	    4'b0110: HEX0 = 7'b0000010;//6
	    4'b0111: HEX0 = 7'b1111000;//7
	    4'b1000: HEX0 = 7'b0000000;//8
	    4'b1001: HEX0 = 7'b0010000;//9
	   4'b1010: HEX0 = 7'b0001000;
		4'b1011: HEX0 = 7'b0000011;
		4'b1100: HEX0 = 7'b1000110;
		4'b1101: HEX0 = 7'b0100001;
		4'b1110: HEX0 = 7'b0000110;
		4'b1111: HEX0 = 7'b0001110;
	endcase 

case (SW[7:4])
	    4'b0000: HEX1 = 7'b1000000;//0
	    4'b0001: HEX1 = 7'b1111001;//1
	    4'b0010: HEX1 = 7'b0100100;//2
	    4'b0011: HEX1 = 7'b0110000;//3
	    4'b0100: HEX1 = 7'b0011001;//4
	    4'b0101: HEX1 = 7'b0010010;//5
	    4'b0110: HEX1 = 7'b0000010;//6
	    4'b0111: HEX1 = 7'b1111000;//7
	    4'b1000: HEX1 = 7'b0000000;//8
	    4'b1001: HEX1 = 7'b0010000;//9
	 4'b1010: HEX1 = 7'b0001000;
		4'b1011: HEX1 = 7'b0000011;
		4'b1100: HEX1 = 7'b1000110;
		4'b1101: HEX1 = 7'b0100001;
		4'b1110: HEX1 = 7'b0000110;
		4'b1111: HEX1 = 7'b0001110;
	endcase
	
case (LEDR[3:0])
	    4'b0000: HEX2 = 7'b1000000;//0
	    4'b0001: HEX2 = 7'b1111001;//1
	    4'b0010: HEX2 = 7'b0100100;//2
	    4'b0011: HEX2 = 7'b0110000;//3
	    4'b0100: HEX2 = 7'b0011001;//4
	    4'b0101: HEX2 = 7'b0010010;//5
	    4'b0110: HEX2 = 7'b0000010;//6
	    4'b0111: HEX2 = 7'b1111000;//7
	    4'b1000: HEX2 = 7'b0000000;//8
	    4'b1001: HEX2 = 7'b0010000;//9
	  4'b1010: HEX2 = 7'b0001000;
		4'b1011: HEX2 = 7'b0000011;
		4'b1100: HEX2 = 7'b1000110;
		4'b1101: HEX2 = 7'b0100001;
		4'b1110: HEX2 = 7'b0000110;
		4'b1111: HEX2 = 7'b0001110;
	endcase 
	
case (LEDR[7:4])
	    4'b0000: HEX3 = 7'b1000000;//0
	    4'b0001: HEX3 = 7'b1111001;//1
	    4'b0010: HEX3 = 7'b0100100;//2
	    4'b0011: HEX3 = 7'b0110000;//3
	    4'b0100: HEX3 = 7'b0011001;//4
	    4'b0101: HEX3 = 7'b0010010;//5
	    4'b0110: HEX3 = 7'b0000010;//6
	    4'b0111: HEX3 = 7'b1111000;//7
	    4'b1000: HEX3 = 7'b0000000;//8
	    4'b1001: HEX3 = 7'b0010000;//9
	   4'b1010: HEX3 = 7'b0001000;
		4'b1011: HEX3 = 7'b0000011;
		4'b1100: HEX3 = 7'b1000110;
		4'b1101: HEX3 = 7'b0100001;
		4'b1110: HEX3 = 7'b0000110;
		4'b1111: HEX3 = 7'b0001110;
	endcase 
end 
endmodule 

						